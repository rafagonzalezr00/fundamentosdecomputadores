
Started : "Simulate Behavioral Model".

Determining files marked for global include in the design...
Running fuse...
Command Line: fuse -intstyle ise -incremental -lib secureip -o D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5_isim_beh.exe -prj D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5_beh.prj work.T_p5 {}
Running: C:\Xilinx\14.7\ISE_DS\ISE\bin\nt64\unwrapped\fuse.exe -intstyle ise -incremental -lib secureip -o D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5_isim_beh.exe -prj D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5_beh.prj work.T_p5 
ISim P.20131013 (signature 0x7708f090)
Number of CPUs detected in this system: 12
Turning on mult-threading, number of parallel sub-compilation jobs: 24 
Determining compilation order of HDL files
Parsing VHDL file "D:/practrica5/practica5_rafaelgonzalez_pablosaldana/practica5.vhd" into library work
Parsing VHDL file "D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5.vhd" into library work
Starting static elaboration
Completed static elaboration
Compiling package standard
Compiling package std_logic_1164
Compiling package std_logic_arith
Compiling package std_logic_unsigned
Compiling architecture behavioral of entity practica5 [practica5_default]
Compiling architecture behavior of entity t_p5
Time Resolution for simulation is 1ps.
WARNING:Simulator - Unable to copy libPortabilityNOSH.dll to the simulation executable directory: boost::filesystem::copy_file: El sistema no puede encontrar la ruta especificada, "isim\T_p5_isim_beh.exe.sim\libPortability.dll".
Compiled 7 VHDL Units
Built simulation executable D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5_isim_beh.exe
Fuse Memory Usage: 34496 KB
Fuse CPU Usage: 327 ms
Launching ISim simulation engine GUI...
"D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5_isim_beh.exe" -intstyle ise -gui -tclbatch isim.cmd  -view "D:/practrica5/practica5_rafaelgonzalez_pablosaldana/p5.wcfg" -wdb "D:/practrica5/practica5_rafaelgonzalez_pablosaldana/T_p5_isim_beh.wdb"
ISim simulation engine GUI launched successfully

Process "Simulate Behavioral Model" completed successfully
